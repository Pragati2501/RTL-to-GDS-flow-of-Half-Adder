magic
tech scmos
magscale 1 2
timestamp 1687607595
<< metal1 >>
rect 280 206 286 214
rect 294 206 300 214
rect 308 206 314 214
rect 322 206 328 214
rect 28 136 32 144
rect 96 142 100 144
rect 109 137 124 143
rect 132 137 179 143
rect 269 137 316 143
rect 236 132 244 136
rect 332 132 340 136
rect 172 124 180 128
rect 120 6 126 14
rect 134 6 140 14
rect 148 6 154 14
rect 162 6 168 14
<< m2contact >>
rect 286 206 294 214
rect 300 206 308 214
rect 314 206 322 214
rect 12 136 20 144
rect 124 136 132 144
rect 316 136 324 144
rect 364 136 372 144
rect 60 116 68 124
rect 188 116 196 124
rect 220 116 228 124
rect 236 116 244 124
rect 332 116 340 124
rect 126 6 134 14
rect 140 6 148 14
rect 154 6 162 14
<< metal2 >>
rect 125 144 131 243
rect 365 237 396 243
rect 280 214 328 216
rect 280 206 282 214
rect 294 206 300 214
rect 308 206 314 214
rect 326 206 328 214
rect 280 204 328 206
rect 365 164 371 237
rect 317 144 323 156
rect 13 124 19 136
rect 365 124 371 136
rect 61 84 67 116
rect 237 84 243 116
rect 120 14 168 16
rect 120 6 122 14
rect 134 6 140 14
rect 148 6 154 14
rect 166 6 168 14
rect 120 4 168 6
<< m3contact >>
rect 282 206 286 214
rect 286 206 290 214
rect 300 206 308 214
rect 318 206 322 214
rect 322 206 326 214
rect 396 236 404 244
rect 316 156 324 164
rect 364 156 372 164
rect 12 116 20 124
rect 188 116 196 124
rect 220 116 228 124
rect 332 116 340 124
rect 364 116 372 124
rect 60 76 68 84
rect 236 76 244 84
rect 122 6 126 14
rect 126 6 130 14
rect 140 6 148 14
rect 158 6 162 14
rect 162 6 166 14
<< metal3 >>
rect 394 244 406 246
rect 394 236 396 244
rect 404 236 406 244
rect 394 234 406 236
rect 280 214 328 216
rect 280 206 282 214
rect 290 206 300 214
rect 308 206 318 214
rect 326 206 328 214
rect 280 204 328 206
rect 395 195 405 234
rect 314 165 326 166
rect 362 165 374 166
rect -21 125 -11 165
rect 314 164 374 165
rect 314 156 316 164
rect 324 156 364 164
rect 372 156 374 164
rect 314 155 374 156
rect 314 154 326 155
rect 362 154 374 155
rect 10 125 22 126
rect 186 125 198 126
rect -21 124 198 125
rect -21 116 12 124
rect 20 116 188 124
rect 196 116 198 124
rect -21 115 198 116
rect 10 114 22 115
rect 186 114 198 115
rect 218 125 230 126
rect 330 125 342 126
rect 218 124 342 125
rect 218 116 220 124
rect 228 116 332 124
rect 340 116 342 124
rect 218 115 342 116
rect 218 114 230 115
rect 330 114 342 115
rect 362 125 374 126
rect 395 125 405 165
rect 362 124 405 125
rect 362 116 364 124
rect 372 116 405 124
rect 362 115 405 116
rect 362 114 374 115
rect 58 85 70 86
rect 234 85 246 86
rect 58 84 246 85
rect 58 76 60 84
rect 68 76 236 84
rect 244 76 246 84
rect 58 75 246 76
rect 58 74 70 75
rect 234 74 246 75
rect 120 14 168 16
rect 120 6 122 14
rect 130 6 140 14
rect 148 6 158 14
rect 166 6 168 14
rect 120 4 168 6
use FILL  FILL_0_0_0
timestamp 1687607595
transform 1 0 120 0 -1 210
box -4 -6 20 206
use XOR2X1  XOR2X1_1
timestamp 1687607595
transform -1 0 120 0 -1 210
box -4 -6 116 206
use BUFX2  BUFX2_2
timestamp 1687607595
transform 1 0 232 0 -1 210
box -4 -6 52 206
use FILL  FILL_0_0_2
timestamp 1687607595
transform 1 0 152 0 -1 210
box -4 -6 20 206
use FILL  FILL_0_0_1
timestamp 1687607595
transform 1 0 136 0 -1 210
box -4 -6 20 206
use AND2X2  AND2X2_1
timestamp 1687607595
transform 1 0 168 0 -1 210
box -4 -6 68 206
use BUFX2  BUFX2_1
timestamp 1687607595
transform 1 0 328 0 -1 210
box -4 -6 52 206
use FILL  FILL_0_1_2
timestamp 1687607595
transform 1 0 312 0 -1 210
box -4 -6 20 206
use FILL  FILL_0_1_1
timestamp 1687607595
transform 1 0 296 0 -1 210
box -4 -6 20 206
use FILL  FILL_0_1_0
timestamp 1687607595
transform 1 0 280 0 -1 210
box -4 -6 20 206
<< labels >>
flabel metal3 s -16 160 -16 160 7 FreeSans 16 0 0 0 a
port 0 nsew
flabel metal2 s 128 240 128 240 3 FreeSans 16 90 0 0 b
port 1 nsew
flabel metal3 s 400 200 400 200 3 FreeSans 16 90 0 0 s
port 2 nsew
flabel metal3 s 400 160 400 160 3 FreeSans 16 0 0 0 c
port 3 nsew
<< end >>
