* NGSPICE file created from half_adder.ext - technology: scmos

* Black-box entry subcircuit for FILL abstract view
.subckt FILL gnd vdd
.ends

* Black-box entry subcircuit for XOR2X1 abstract view
.subckt XOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for BUFX2 abstract view
.subckt BUFX2 A gnd Y vdd
.ends

* Black-box entry subcircuit for AND2X2 abstract view
.subckt AND2X2 A B gnd Y vdd
.ends

.subckt half_adder a b s c
XFILL_0_0_0 BUFX2_2/gnd BUFX2_2/vdd FILL
XFILL_0_0_1 BUFX2_2/gnd BUFX2_2/vdd FILL
XFILL_0_0_2 BUFX2_2/gnd BUFX2_2/vdd FILL
XXOR2X1_1 b a BUFX2_2/gnd BUFX2_2/A BUFX2_2/vdd XOR2X1
XBUFX2_1 BUFX2_1/A BUFX2_2/gnd c BUFX2_2/vdd BUFX2
XBUFX2_2 BUFX2_2/A BUFX2_2/gnd s BUFX2_2/vdd BUFX2
XFILL_0_1_0 BUFX2_2/gnd BUFX2_2/vdd FILL
XFILL_0_1_1 BUFX2_2/gnd BUFX2_2/vdd FILL
XFILL_0_1_2 BUFX2_2/gnd BUFX2_2/vdd FILL
XAND2X2_1 b a BUFX2_2/gnd BUFX2_1/A BUFX2_2/vdd AND2X2
.ends

