VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO half_adder
  CLASS BLOCK ;
  FOREIGN half_adder ;
  ORIGIN 3.150 -0.600 ;
  SIZE 64.050 BY 36.300 ;
  PIN a
    PORT
      LAYER metal1 ;
        RECT 1.800 20.400 3.000 21.600 ;
        RECT 28.200 17.400 29.400 18.600 ;
      LAYER metal2 ;
        RECT 1.800 20.400 3.000 21.600 ;
        RECT 1.950 18.600 2.850 20.400 ;
        RECT 1.800 17.400 3.000 18.600 ;
        RECT 28.200 17.400 29.400 18.600 ;
      LAYER metal3 ;
        RECT -3.150 18.750 -1.650 24.750 ;
        RECT 1.500 18.750 3.300 18.900 ;
        RECT 27.900 18.750 29.700 18.900 ;
        RECT -3.150 17.250 29.700 18.750 ;
        RECT 1.500 17.100 3.300 17.250 ;
        RECT 27.900 17.100 29.700 17.250 ;
    END
  END a
  PIN b
    PORT
      LAYER metal1 ;
        RECT 16.200 21.450 17.400 21.600 ;
        RECT 18.600 21.450 19.800 21.600 ;
        RECT 25.800 21.450 27.000 21.600 ;
        RECT 16.200 20.550 27.000 21.450 ;
        RECT 16.200 20.400 17.400 20.550 ;
        RECT 18.600 20.400 19.800 20.550 ;
        RECT 25.800 20.400 27.000 20.550 ;
      LAYER metal2 ;
        RECT 18.750 21.600 19.650 36.450 ;
        RECT 18.600 20.400 19.800 21.600 ;
    END
  END b
  PIN s
    PORT
      LAYER metal1 ;
        RECT 40.200 21.450 41.400 21.600 ;
        RECT 47.400 21.450 48.600 21.600 ;
        RECT 40.200 20.550 48.600 21.450 ;
        RECT 40.200 20.400 41.400 20.550 ;
        RECT 47.400 20.400 48.600 20.550 ;
      LAYER metal2 ;
        RECT 59.400 36.450 60.600 36.600 ;
        RECT 54.750 35.550 60.600 36.450 ;
        RECT 54.750 24.600 55.650 35.550 ;
        RECT 59.400 35.400 60.600 35.550 ;
        RECT 47.400 23.400 48.600 24.600 ;
        RECT 54.600 23.400 55.800 24.600 ;
        RECT 47.550 21.600 48.450 23.400 ;
        RECT 47.400 20.400 48.600 21.600 ;
      LAYER metal3 ;
        RECT 59.100 35.100 60.900 36.900 ;
        RECT 59.250 29.250 60.750 35.100 ;
        RECT 47.100 24.750 48.900 24.900 ;
        RECT 54.300 24.750 56.100 24.900 ;
        RECT 47.100 23.250 56.100 24.750 ;
        RECT 47.100 23.100 48.900 23.250 ;
        RECT 54.300 23.100 56.100 23.250 ;
    END
  END s
  PIN c
    PORT
      LAYER metal1 ;
        RECT 54.600 20.400 55.800 21.600 ;
      LAYER metal2 ;
        RECT 54.600 20.400 55.800 21.600 ;
        RECT 54.750 18.600 55.650 20.400 ;
        RECT 54.600 17.400 55.800 18.600 ;
      LAYER metal3 ;
        RECT 54.300 18.750 56.100 18.900 ;
        RECT 59.250 18.750 60.750 24.750 ;
        RECT 54.300 17.250 60.750 18.750 ;
        RECT 54.300 17.100 56.100 17.250 ;
    END
  END c
  OBS
      LAYER metal1 ;
        RECT 0.600 30.600 57.000 32.400 ;
        RECT 1.800 23.700 3.000 29.700 ;
        RECT 4.200 24.600 5.700 29.700 ;
        RECT 8.400 24.300 10.800 29.700 ;
        RECT 13.500 24.600 15.000 29.700 ;
        RECT 1.800 22.800 5.400 23.700 ;
        RECT 4.200 22.500 5.400 22.800 ;
        RECT 6.300 22.200 7.500 23.400 ;
        RECT 6.300 21.600 7.200 22.200 ;
        RECT 3.900 20.400 4.800 21.600 ;
        RECT 6.000 20.400 7.200 21.600 ;
        RECT 8.400 21.300 9.300 24.300 ;
        RECT 16.200 23.700 17.400 29.700 ;
        RECT 25.800 23.700 27.000 29.700 ;
        RECT 29.700 24.000 30.900 29.700 ;
        RECT 32.100 25.200 33.300 29.700 ;
        RECT 32.100 23.700 34.200 25.200 ;
        RECT 10.200 22.200 12.600 23.400 ;
        RECT 13.500 22.800 17.400 23.700 ;
        RECT 26.100 23.400 27.000 23.700 ;
        RECT 26.100 22.800 28.800 23.400 ;
        RECT 13.500 22.500 14.700 22.800 ;
        RECT 26.100 22.500 32.400 22.800 ;
        RECT 27.900 21.900 32.400 22.500 ;
        RECT 31.200 21.600 32.400 21.900 ;
        RECT 14.400 21.300 15.300 21.600 ;
        RECT 8.400 20.400 9.900 21.300 ;
        RECT 14.100 21.000 15.300 21.300 ;
        RECT 9.000 19.500 9.900 20.400 ;
        RECT 10.800 20.400 15.300 21.000 ;
        RECT 28.800 20.700 30.000 21.000 ;
        RECT 10.800 20.100 15.000 20.400 ;
        RECT 10.800 19.800 12.000 20.100 ;
        RECT 28.500 19.800 30.000 20.700 ;
        RECT 28.500 19.500 29.400 19.800 ;
        RECT 25.800 18.600 27.000 19.500 ;
        RECT 9.000 17.400 10.200 18.600 ;
        RECT 12.900 18.300 14.100 18.600 ;
        RECT 11.700 17.400 14.100 18.300 ;
        RECT 11.700 17.100 12.900 17.400 ;
        RECT 31.200 16.500 32.100 21.600 ;
        RECT 33.300 19.500 34.200 23.700 ;
        RECT 35.400 22.800 36.600 29.700 ;
        RECT 37.800 23.700 39.000 29.700 ;
        RECT 35.400 21.900 38.700 22.800 ;
        RECT 40.200 22.500 41.400 29.700 ;
        RECT 49.800 22.800 51.000 29.700 ;
        RECT 52.200 23.700 53.400 29.700 ;
        RECT 49.800 21.900 53.100 22.800 ;
        RECT 54.600 22.500 55.800 29.700 ;
        RECT 35.400 19.500 36.600 20.400 ;
        RECT 33.000 17.400 34.200 18.600 ;
        RECT 35.400 17.400 36.600 18.600 ;
        RECT 37.800 17.400 38.700 21.900 ;
        RECT 49.800 19.500 51.000 20.400 ;
        RECT 40.200 18.600 41.400 19.500 ;
        RECT 9.000 15.300 9.900 16.500 ;
        RECT 28.500 15.600 32.100 16.500 ;
        RECT 1.800 14.400 5.400 15.300 ;
        RECT 1.800 3.300 3.000 14.400 ;
        RECT 4.200 14.100 5.400 14.400 ;
        RECT 4.200 3.300 5.700 13.200 ;
        RECT 8.400 3.300 10.800 15.300 ;
        RECT 13.500 14.400 17.400 15.300 ;
        RECT 13.500 14.100 14.700 14.400 ;
        RECT 13.500 3.300 15.000 13.200 ;
        RECT 16.200 3.300 17.400 14.400 ;
        RECT 28.500 9.300 29.400 15.600 ;
        RECT 33.300 15.300 34.200 16.500 ;
        RECT 37.800 16.200 39.600 17.400 ;
        RECT 37.800 15.300 38.700 16.200 ;
        RECT 40.500 15.300 41.400 18.600 ;
        RECT 49.800 17.400 51.000 18.600 ;
        RECT 52.200 17.400 53.100 21.900 ;
        RECT 54.600 18.600 55.800 19.500 ;
        RECT 52.200 16.200 54.000 17.400 ;
        RECT 52.200 15.300 53.100 16.200 ;
        RECT 54.900 15.300 55.800 18.600 ;
        RECT 25.800 3.300 27.000 9.300 ;
        RECT 28.200 3.300 29.400 9.300 ;
        RECT 30.600 3.300 31.800 14.700 ;
        RECT 33.000 3.300 34.200 15.300 ;
        RECT 35.400 14.400 38.700 15.300 ;
        RECT 35.400 3.300 36.600 14.400 ;
        RECT 37.800 3.300 39.000 13.500 ;
        RECT 40.200 3.300 41.400 15.300 ;
        RECT 49.800 14.400 53.100 15.300 ;
        RECT 49.800 3.300 51.000 14.400 ;
        RECT 52.200 3.300 53.400 13.500 ;
        RECT 54.600 3.300 55.800 15.300 ;
        RECT 0.600 0.600 57.000 2.400 ;
      LAYER via1 ;
        RECT 42.900 30.900 44.100 32.100 ;
        RECT 45.000 30.900 46.200 32.100 ;
        RECT 47.100 30.900 48.300 32.100 ;
        RECT 11.400 22.200 12.600 23.400 ;
        RECT 18.900 0.900 20.100 2.100 ;
        RECT 21.000 0.900 22.200 2.100 ;
        RECT 23.100 0.900 24.300 2.100 ;
      LAYER metal2 ;
        RECT 42.000 30.600 49.200 32.400 ;
        RECT 4.200 22.500 5.400 23.700 ;
        RECT 13.500 23.400 14.700 23.700 ;
        RECT 6.300 22.500 14.700 23.400 ;
        RECT 4.200 21.300 5.100 22.500 ;
        RECT 6.300 22.200 7.500 22.500 ;
        RECT 11.400 22.200 12.600 22.500 ;
        RECT 4.200 20.400 12.600 21.300 ;
        RECT 4.200 15.300 5.100 20.400 ;
        RECT 9.000 17.400 10.200 18.600 ;
        RECT 11.700 18.300 12.600 20.400 ;
        RECT 4.200 14.100 5.400 15.300 ;
        RECT 9.150 12.600 10.050 17.400 ;
        RECT 11.700 17.100 12.900 18.300 ;
        RECT 13.800 15.300 14.700 22.500 ;
        RECT 33.000 17.400 34.200 18.600 ;
        RECT 35.400 17.400 36.600 18.600 ;
        RECT 49.800 17.400 51.000 18.600 ;
        RECT 13.500 14.100 14.700 15.300 ;
        RECT 35.550 12.600 36.450 17.400 ;
        RECT 9.000 11.400 10.200 12.600 ;
        RECT 35.400 11.400 36.600 12.600 ;
        RECT 18.000 0.600 25.200 2.400 ;
      LAYER via2 ;
        RECT 42.300 30.900 43.500 32.100 ;
        RECT 45.000 30.900 46.200 32.100 ;
        RECT 47.700 30.900 48.900 32.100 ;
        RECT 18.300 0.900 19.500 2.100 ;
        RECT 21.000 0.900 22.200 2.100 ;
        RECT 23.700 0.900 24.900 2.100 ;
      LAYER metal3 ;
        RECT 42.000 30.600 49.200 32.400 ;
        RECT 32.700 18.750 34.500 18.900 ;
        RECT 49.500 18.750 51.300 18.900 ;
        RECT 32.700 17.250 51.300 18.750 ;
        RECT 32.700 17.100 34.500 17.250 ;
        RECT 49.500 17.100 51.300 17.250 ;
        RECT 8.700 12.750 10.500 12.900 ;
        RECT 35.100 12.750 36.900 12.900 ;
        RECT 8.700 11.250 36.900 12.750 ;
        RECT 8.700 11.100 10.500 11.250 ;
        RECT 35.100 11.100 36.900 11.250 ;
        RECT 18.000 0.600 25.200 2.400 ;
  END
END half_adder
END LIBRARY

